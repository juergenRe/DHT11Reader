----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/01/2020 10:26:36 AM
-- Design Name: 
-- Module Name: DHT11Control_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DHT11Control_tb is
end DHT11Control_tb;

architecture Behavioral of DHT11Control_tb is
   -- Clock period definitions
constant clk_period:    time := 10 ns;

   --internal signals
signal clk:             std_logic := '0';
signal reset:           std_logic := '0';

-- inputs to DHT11Reader block
constant NDIV:          integer := 99;

signal outT:           std_logic_vector(15 downto 0);      -- temperature
signal outH:           std_logic_vector(15 downto 0);      -- humidity
signal outStatus:      std_logic_vector(1 downto 0);       -- status: [1]: sample available; [0]: error
signal rdy:            std_logic;                          -- component ready to receive new settings
signal dhtOutSig:      std_logic;                          -- driver line to DHT11

signal trg:            std_logic := '0';                   -- new settings trigger
signal dhtInSig:       std_logic := '1';                   -- input line towards simulated DHT11

-----------------------------------
-- dht11 simulation signals
--
constant NDATABIT:      integer := 40;
signal txData:          std_logic_vector(NDATABIT-1 downto 0) := (others => '0');

-- timing constants: base timing, can be streteched by MULT
-- times are nominal times
constant MULT:          integer := 5;
constant TSTRTIN:       time := 10us;               -- min time to detect a trigger
constant TWAKE:         time := 30us;               -- wake up 20..40us
constant TSTRTL:        time := 80us;               -- duration of start bit low of DHT
constant TSTRTH:        time := 80us;               -- duration of start bit high
constant TBITL:         time := 50us;               -- duration of bit low time
constant TBITH0:        time := 27us;               -- duration of bit high when transmitting '0'
constant TBITH1:        time := 70us;               -- duration of bit high when transmitting '1'
constant TEXCESSTIME:   time := 17ms;               -- excessive hold of one state

constant TVAR_WAKE_MN:  time := 10us;               -- variation to get minimum time 
constant TVAR_WAKE_MX:  time := 10us;               -- variation to get maximum time 
constant TVAR_STRT_MN:  time := 20us;               -- variation to get minimum time 
constant TVAR_STRT_MX:  time := 20us;               -- variation to get maximum time 
constant TVAR_BITL_MN:  time := 10us;               -- variation to get minimum time 
constant TVAR_BITL_MX:  time := 10us;               -- variation to get maximum time 
constant TVAR_BITH0_MN: time :=  7us;               -- variation to get minimum time 
constant TVAR_BITH0_MX: time := 13us;               -- variation to get maximum time 
constant TVAR_BITH1_MN: time := 10us;               -- variation to get minimum time 
constant TVAR_BITH1_MX: time := 10us;               -- variation to get maximum time 

constant TD_ERROR:      time :=  1us;               -- additaional time increment to get out of good window

signal t_trigin:        time;                   -- min external start bit
signal t_wakeup:        time;
signal t_startL:        time;
signal t_startH:        time;
signal t_bitL:          time;
signal t_bitH0:         time;
signal t_bitH1:         time;

-- Test Data definiton
constant NB_TIMES:      natural := 7;
type t_timing_ary is array (natural range <>) of time;
type t_testdata is record
      timings   : t_timing_ary(0 to NB_TIMES-1);	-- timing array
	  data	    : std_logic_vector(31 downto 0); 	-- data to transmit
	  expectRes	: boolean;						    -- expected result
	  expectSC  : boolean;                          -- expected short circuit detection
	  desc      : string(1 to 40);                  -- description string
end record;
type t_test_ary is array (natural range <>) of t_testdata;

  ------------------------------------------------------------------------------
  -- Stimulus data
  ------------------------------------------------------------------------------
  -- The following constant holds the stimulus for the testbench. It is
  -- an ordered array of timings and data to transmit.
  ------------------------------------------------------------------------------
constant test_data : t_test_ary := (
    0       => (            -- good timing
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => false,
      expectSC => false,
      desc      => "<0> Good timings A                      "),
    1       => (            -- good timing
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"00000000",
      expectRes => false,
      expectSC => false,
      desc      => "<1> Good timings B                      "),
    2       => (            -- good timing
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"FFFFFFFF",
      expectRes => false,
      expectSC => false,
      desc      => "<2> Good timings C                      "),
    3       => (            -- wake up too long
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE + TVAR_WAKE_MX + TD_ERROR,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<3> Wake up too long                    "),
    4       => (            -- Start bit "0" DHT too short
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL - TVAR_STRT_MN - TD_ERROR,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<4> Start bit DHT too short             "),
    5       => (            -- Start bit "0" DHT too long
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL + TVAR_STRT_MX + TD_ERROR,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<5> Start bit DHT too long              "),
    6       => (            -- Start bit "1" DHT too short
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH - TVAR_STRT_MN - TD_ERROR,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<6> Start bit DHT High too short        "),
    7       => (            -- Start bit "1" DHT too long
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH + TVAR_STRT_MX + TD_ERROR,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<7> Start bit DHT High too long         "),
    8       => (            -- TXLow phase too short
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,
                     4 => TBITL - TVAR_BITL_MN - TD_ERROR,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<8> TX Bit low too short                "),
    9       => (            -- TXLow phase too long
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL + TVAR_BITL_MX + TD_ERROR,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<9> TX Bit low too long                 "),
    10      => (            -- TXHigh phase too short (less than '0' bit length)
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,
                     4 => TBITL,  
                     5 => TBITH0 - TVAR_BITH0_MN - TD_ERROR,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<10> TX Bit High too short for '0'      "),
      --           "0123456789012345678901234567890123456789"
    11      => (            -- TXHigh phase too long for '0'
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0 + TVAR_BITH0_MX + TD_ERROR,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<11> TX Bit High too long for '0'       "),
      --           "0123456789012345678901234567890123456789"
    12      => (            -- TXHigh phase too short for '1'
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1 - TVAR_BITH1_MN - TD_ERROR),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<12> TX Bit High too short for '1'      "),
      --           "0123456789012345678901234567890123456789"
    13      => (            -- TXHigh phase too long for '1'
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1 + TVAR_BITH1_MX + TD_ERROR),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<13> TX Bit High too long for '1'       "),
    14      => (            -- repeat good timing to check if status is reset correctly
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => false,
      expectSC => false,
      desc      => "<14> Good timings A (repeat)            "),
    15      => (            -- excessive start bit low --> counter overflow
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TEXCESSTIME,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => true,
      desc      => "<15> Excess start bit L                 "),
    16      => (            -- excessive start bit high --> counter overflow
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TEXCESSTIME,  
                     4 => TBITL,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<16> Excess start bit H                 "),
    17      => (            -- excessive Tx bit high --> counter overflow
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TEXCESSTIME,  
                     5 => TBITH0,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => true,
      desc      => "<17> Excess Tx bit L                    "),
    18      => (            -- excessive Tx bit low --> counter overflow
      timings   => ( 0 => TSTRTIN,
                     1 => TWAKE,
                     2 => TSTRTL,  
                     3 => TSTRTH,  
                     4 => TBITL,  
                     5 => TEXCESSTIME,  
                     6 => TBITH1),
      data      => x"5577AA33",
      expectRes => true,
      expectSC => false,
      desc      => "<18> Excess Tx bit H                    ")
      --           "0123456789012345678901234567890123456789"
      ); 

type t_testState is (stPowOn, stIdle, stTestSetUp, stTestStart, stTestRun, stTestEnd);
signal testStateReg:    t_testState;
signal testStateNxt:    t_testState;
signal startTest:       std_logic;
signal testDone:        std_logic;
signal testCnt:         unsigned(4 downto 0);       -- holds the current test index

----------------------------------------------------------------
signal expectResult:boolean;

----------------------------------------
component DHT11Control
    generic (
        NDIV:           integer := 99;                          -- 1us ticks @ 100MHz clock
        POWONDLY:       boolean := false                        -- enable simulation timings or real timings
    );
    port (
        clk:            in std_logic;
        reset:          in std_logic;
        cntTick:        out std_logic;                          -- counter tick
        outT:           out std_logic_vector(15 downto 0);      -- temperature out
        outH:           out std_logic_vector(15 downto 0);      -- humidity out
        outStatus:      out std_logic_vector(1 downto 0);       -- status out: [1]: sample available; [0]: error
        trg:            in std_logic;                           -- new settings trigger
        rdy:            out std_logic;                          -- component ready to receive new settings
        dhtInSig:       in std_logic;                           -- input line from DHT11
        dhtOutSig:      out std_logic                           -- output line to DHT11
     );
end component;

component DHT11DeviceSimulation is
    generic (
        NDATABIT:      integer := 40
    );
    port (
        clk:            in std_logic;
        reset:          in std_logic;
        dhtInSig:       out std_logic;                          -- input line from DHT11
        dhtOutSig:      in std_logic;                           -- output line to DHT11
        -- configuration inputs for device
        t_trigin:       in time;
        t_wakeup:       in time;
        t_startL:       in time;
        t_startH:       in time;
        t_bitL:         in time;
        t_bitH0:        in time;
        t_bitH1:        in time;
        txData:         in std_logic_vector(NDATABIT-1 downto 0)
     );
end component;

procedure wrOut (arg : in string := "") is
begin
  std.textio.write(std.textio.output, arg & LF);
end procedure wrOut;

begin
    uut: DHT11Control
        generic map(
            NDIV        => NDIV,  
            POWONDLY    => false
        )
        port map (
            clk         => clk,     
            reset       => reset,
            cntTick     => open,
            outT        => outT,
            outH        => outH,
            outStatus   => outStatus,
            trg         => trg,
            rdy         => rdy,
            dhtInSig    => dhtInSig,
            dhtOutSig   => dhtOutSig
         );

    dht11_dvc: DHT11DeviceSimulation
        generic map (     
            NDATABIT    => NDATABIT
        )          
        port map (        
            clk         => clk,
            reset       => reset,
            dhtInSig    => dhtInSig,
            dhtOutSig   => dhtOutSig,
            t_trigin    => t_trigin, 
            t_wakeup    => t_wakeup,
            t_startL    => t_startL,
            t_startH    => t_startH,
            t_bitL      => t_bitL, 
            t_bitH0     => t_bitH0,
            t_bitH1     => t_bitH1,  
            txData      => txData    
         );           	
    
 -------------------------------------------------------------------   
 -- Clock process definitions                                            
    clk_process :process
	begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
	end process;

   -------------------------------------------------------------------
   -- Stimulus process
    stim_proc: process
    begin
        -- check behaviour when no reset is given
        startTest <= '0';
        wait for 200 ns;
        reset <= '1';
        wait for 100ns;
        reset <= '0';
		wait until rdy = '1';
		wait for 200ns;
		wait until rising_edge(clk);
		--wait until testDone = '1';
		startTest <= '1';
		wait until rising_edge(clk);
		wait until testDone = '0';
		wait until rising_edge(clk);
		startTest <= '0';
		wait until testDone = '1';
		
		wait for 100ns;
		assert false report "Simulation done" severity failure;
	end process;
	

----------------------------------------------------------------------------------
-- traverse through test sets triggered by trg signal
    dht11_test_pattern_reg: process(clk, reset)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                testStateReg <= stPowOn;
            else
                testStateReg <= testStateNxt;
            end if;
        end if;
    end process dht11_test_pattern_reg;
    
    testDone <= '1' when (testStateReg = stIdle) else '0';

    dht11_test_pattern_nxt: process(testStateReg, startTest, rdy)
        variable actIdx:    integer := 0;
        variable dataVal:   std_logic_vector(31 downto 0);
        variable er:        boolean;
        variable sc:        boolean;
        variable desc:      string(1 to 40);
        variable res:       integer;
        variable stat:      boolean;
        variable statsc:    boolean;
        
        function calc_crc ( data : in std_logic_vector) return std_logic_vector is
            variable crc: std_logic_vector(7 downto 0);
		begin
		    crc := data(31 downto 24) + data(23 downto 16) + data(15 downto 8) + data(7 downto 0);
		    return crc;
		end;
        procedure getActData(idx: in natural; dx: out std_logic_vector; expectResult: out boolean; expectSC: out boolean; desc: out string) is
        begin
            dx := test_data(idx).data;
            t_trigin <= test_data(idx).timings(0);
            t_wakeup <= test_data(idx).timings(1);
            t_startL <= test_data(idx).timings(2);
            t_startH <= test_data(idx).timings(3);
            t_bitL  <= test_data(idx).timings(4);
            t_bitH0 <= test_data(idx).timings(5);
            t_bitH1 <= test_data(idx).timings(6);
            expectResult := test_data(idx).expectRes;
            expectSC := test_data(idx).expectSC;
            desc := test_data(idx).desc;
        end;
    begin
        case testStateReg is
            when stPowOn =>
                testStateNxt <= stIdle;
                testCnt <= (others => '0');
            when stIdle =>
                actIdx := 0;
                if startTest = '1' and rdy = '1' then
                    testStateNxt <= stTestSetUp;
                end if;
            when stTestSetUp =>
                testCnt <= TO_UNSIGNED(actIdx, 5);
                getActData(actIdx, dataVal, er, sc, desc);
                txData <= dataVal & calc_crc(dataVal);
                wrOut("---------------------------------------------");
                wrOut("Start Test: " & desc);
                testStateNxt <= stTestStart;
            when stTestStart =>
                trg <= '1';
                if rdy = '0' then
                    testStateNxt <= stTestRun;
                    trg <= '0';
                end if;
            when stTestRun => 
                -- executing reception, wait till finished
                if rdy = '1' then
                    res := conv_integer(outH & outT);
                    stat := (outStatus(0) = '1');
                    statsc := (outStatus(1) = '1');
                    assert not (er xor stat)
                        report "Expected status unequal expect=" & boolean'image(er) & " => measured=" & boolean'image(stat) severity error;
                        
                    assert not (sc xor statsc)
                        report "Expected short circuit status unequal: expect=" & boolean'image(sc) & " => measured=" & boolean'image(statsc) severity error;
                        
                    if not stat then
                        assert res = conv_integer(dataVal)
                            report "Expected data values unequal data=" & integer'image(conv_integer(dataVal)) & " => outH/T: " & integer'image(res) severity error;
                    end if;

                    testStateNxt <= stTestSetUp;
                    actIdx := actIdx + 1;
                    if actIdx = test_data'length then
                        testStateNxt <= stTestEnd;
                    end if;
                end if;
            when stTestEnd =>
                wrOut("---------------------------------------------");
                wrOut("Test done");
                testStateNxt <= stIdle; 
        end case;
    end process dht11_test_pattern_nxt;
    
end Behavioral;
  
    
   
   
    
   
   
